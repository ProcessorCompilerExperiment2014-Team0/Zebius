library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package zebius is

  subtype reg_data is unsigned(31 downto 0);

end zebius;

